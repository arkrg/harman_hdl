module env_test(
	input a, b,
	output c
);

// an and-gate for testing this simulation enviroment

	assign c = a & b;
endmodule
